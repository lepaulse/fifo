module fifo #(parameter 
                BUFFER_SIZE = 128, // From 1 to 127 values  
                DATA_WIDTH = 32,
                ADDRESS_WIDTH = clogb2(BUFFER_SIZE)
             )
    (
    // Data in interface
    input wire rst_in_n,
    input wire clock_in,
    input wire [DATA_WIDTH-1:0] data_in,
    input wire data_in_valid,
    output wire data_in_full,

    // Data out interface
    input wire rst_out_n,
    input wire clock_out,
    output wire [DATA_WIDTH-1:0] data_out,
    output wire data_out_valid,
    input wire data_out_ack
    );


    reg [DATA_WIDTH-1:0] Buffer[BUFFER_SIZE-1:0];
    reg [DATA_WIDTH-1:0] BufferData = {DATA_WIDTH{1'b0}};

    reg [ADDRESS_WIDTH:0] WritePointer2Read, ReadPointer2Write;


    wire [ADDRESS_WIDTH-1:0] WriteAddress, ReadAddress; // Binary memory address 
    reg [ADDRESS_WIDTH:0] WritePointer, ReadPointer;   // Gray coded Pointers for syncronizing across clock domains


    wire DataInFull;
    assign data_in_full = DataInFull;

    assign WriteAddress = 7'b0000001;
    assign ReadAddress = 7'b0000001;




    // Block ram buffer
    // See XilinxSimpleDualPort1ClockBlockRamExample.v for detailed documentation
    generate
        integer ram_index;
        initial
            for (ram_index = 0; ram_index < BUFFER_SIZE; ram_index = ram_index + 1)
                Buffer[ram_index] = {DATA_WIDTH{1'b0}};
    endgenerate

    always @(posedge clock_in) begin
        if (data_in_valid && !DataInFull)
            Buffer[WriteAddress] <= data_in;
        //if (data_out_valid)
        //BufferData <= Buffer[0];
    end

    //TODO: check ram type generated by adding/remving BufferData register:
    assign data_out = Buffer[ReadAddress];
    //assign data_out = BufferData;

    function integer clogb2;
        input integer depth;
              for (clogb2=0; depth>0; clogb2=clogb2+1)
                    depth = depth >> 1;
    endfunction

    //TEMP DEV LOGIC
    assign DataInFull = 1'b0;

endmodule